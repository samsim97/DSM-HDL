`timescale 1ns/1ps

module tb_top_dsm_dac_order_1;

  parameter integer DATA_WIDTH = 16;
  localparam integer NUM_SAMPLES = 100;
  localparam integer OSR = 64;

  reg r_clk = 0;
  reg r_rst_n = 0;
  reg r_sample = 1;
  reg signed [DATA_WIDTH-1:0] r_data_in = 0;
  wire w_bit_out;

  reg signed [DATA_WIDTH-1:0] r_input_signal [0:NUM_SAMPLES-1];

  initial begin
    // 300 samples test
    r_input_signal[0] = 16'b0000000000000000;
    r_input_signal[1] = 16'b0000000100010010; 
    r_input_signal[2] = 16'b0000001000100100; 
    r_input_signal[3] = 16'b0000001100110110; 
    r_input_signal[4] = 16'b0000010001001000; 
    r_input_signal[5] = 16'b0000010101011010; 
    r_input_signal[6] = 16'b0000011001101010; 
    r_input_signal[7] = 16'b0000011101111010; 
    r_input_signal[8] = 16'b0000100010001001; 
    r_input_signal[9] = 16'b0000100110010111; 
    r_input_signal[10] = 16'b0000101010100101;
    r_input_signal[11] = 16'b0000101110110000;
    r_input_signal[12] = 16'b0000110010111011;
    r_input_signal[13] = 16'b0000110111000100;
    r_input_signal[14] = 16'b0000111011001100;
    r_input_signal[15] = 16'b0000111111010010;
    r_input_signal[16] = 16'b0001000011010110;
    r_input_signal[17] = 16'b0001000111011000;
    r_input_signal[18] = 16'b0001001011011000;
    r_input_signal[19] = 16'b0001001111010111;
    r_input_signal[20] = 16'b0001010011010011;
    r_input_signal[21] = 16'b0001010111001100;
    r_input_signal[22] = 16'b0001011011000011;
    r_input_signal[23] = 16'b0001011110111000;
    r_input_signal[24] = 16'b0001100010101010;
    r_input_signal[25] = 16'b0001100110011001;
    r_input_signal[26] = 16'b0001101010000101;
    r_input_signal[27] = 16'b0001101101101110;
    r_input_signal[28] = 16'b0001110001010101;
    r_input_signal[29] = 16'b0001110100111000;
    r_input_signal[30] = 16'b0001111000010111;
    r_input_signal[31] = 16'b0001111011110100;
    r_input_signal[32] = 16'b0001111111001101;
    r_input_signal[33] = 16'b0010000010100010;
    r_input_signal[34] = 16'b0010000101110100;
    r_input_signal[35] = 16'b0010001001000010;
    r_input_signal[36] = 16'b0010001100001100;
    r_input_signal[37] = 16'b0010001111010010;
    r_input_signal[38] = 16'b0010010010010100;
    r_input_signal[39] = 16'b0010010101010010;
    r_input_signal[40] = 16'b0010011000001100;
    r_input_signal[41] = 16'b0010011011000001;
    r_input_signal[42] = 16'b0010011101110010;
    r_input_signal[43] = 16'b0010100000011111;
    r_input_signal[44] = 16'b0010100011000111;
    r_input_signal[45] = 16'b0010100101101011;
    r_input_signal[46] = 16'b0010101000001010;
    r_input_signal[47] = 16'b0010101010100100;
    r_input_signal[48] = 16'b0010101100111010;
    r_input_signal[49] = 16'b0010101111001011;
    r_input_signal[50] = 16'b0010110001010110;
    r_input_signal[51] = 16'b0010110011011101;
    r_input_signal[52] = 16'b0010110101011111;
    r_input_signal[53] = 16'b0010110111011011;
    r_input_signal[54] = 16'b0010111001010011;
    r_input_signal[55] = 16'b0010111011000101;
    r_input_signal[56] = 16'b0010111100110010;
    r_input_signal[57] = 16'b0010111110011010;
    r_input_signal[58] = 16'b0010111111111100;
    r_input_signal[59] = 16'b0011000001011001;
    r_input_signal[60] = 16'b0011000010110001;
    r_input_signal[61] = 16'b0011000100000011;
    r_input_signal[62] = 16'b0011000101001111;
    r_input_signal[63] = 16'b0011000110010111;
    r_input_signal[64] = 16'b0011000111011000;
    r_input_signal[65] = 16'b0011001000010100;
    r_input_signal[66] = 16'b0011001001001010;
    r_input_signal[67] = 16'b0011001001111011;
    r_input_signal[68] = 16'b0011001010100110;
    r_input_signal[69] = 16'b0011001011001011;
    r_input_signal[70] = 16'b0011001011101010;
    r_input_signal[71] = 16'b0011001100000100;
    r_input_signal[72] = 16'b0011001100011000;
    r_input_signal[73] = 16'b0011001100100111;
    r_input_signal[74] = 16'b0011001100101111;
    r_input_signal[75] = 16'b0011001100110010;
    r_input_signal[76] = 16'b0011001100101111;
    r_input_signal[77] = 16'b0011001100100111;
    r_input_signal[78] = 16'b0011001100011000;
    r_input_signal[79] = 16'b0011001100000100;
    r_input_signal[80] = 16'b0011001011101010;
    r_input_signal[81] = 16'b0011001011001011;
    r_input_signal[82] = 16'b0011001010100110;
    r_input_signal[83] = 16'b0011001001111011;
    r_input_signal[84] = 16'b0011001001001010;
    r_input_signal[85] = 16'b0011001000010100;
    r_input_signal[86] = 16'b0011000111011000;
    r_input_signal[87] = 16'b0011000110010111;
    r_input_signal[88] = 16'b0011000101001111;
    r_input_signal[89] = 16'b0011000100000011;
    r_input_signal[90] = 16'b0011000010110001;
    r_input_signal[91] = 16'b0011000001011001;
    r_input_signal[92] = 16'b0010111111111100;
    r_input_signal[93] = 16'b0010111110011010;
    r_input_signal[94] = 16'b0010111100110010;
    r_input_signal[95] = 16'b0010111011000101;
    r_input_signal[96] = 16'b0010111001010011;
    r_input_signal[97] = 16'b0010110111011011;
    r_input_signal[98] = 16'b0010110101011111;
    r_input_signal[99] = 16'b0010110011011101;
    r_input_signal[100] = 16'b0010110001010110;
    r_input_signal[101] = 16'b0010101111001011;
    r_input_signal[102] = 16'b0010101100111010;
    r_input_signal[103] = 16'b0010101010100100;
    r_input_signal[104] = 16'b0010101000001010;
    r_input_signal[105] = 16'b0010100101101011;
    r_input_signal[106] = 16'b0010100011000111;
    r_input_signal[107] = 16'b0010100000011111;
    r_input_signal[108] = 16'b0010011101110010;
    r_input_signal[109] = 16'b0010011011000001;
    r_input_signal[110] = 16'b0010011000001100;
    r_input_signal[111] = 16'b0010010101010010;
    r_input_signal[112] = 16'b0010010010010100;
    r_input_signal[113] = 16'b0010001111010010;
    r_input_signal[114] = 16'b0010001100001100;
    r_input_signal[115] = 16'b0010001001000010;
    r_input_signal[116] = 16'b0010000101110100;
    r_input_signal[117] = 16'b0010000010100010;
    r_input_signal[118] = 16'b0001111111001101;
    r_input_signal[119] = 16'b0001111011110100;
    r_input_signal[120] = 16'b0001111000010111;
    r_input_signal[121] = 16'b0001110100111000;
    r_input_signal[122] = 16'b0001110001010101;
    r_input_signal[123] = 16'b0001101101101110;
    r_input_signal[124] = 16'b0001101010000101;
    r_input_signal[125] = 16'b0001100110011001;
    r_input_signal[126] = 16'b0001100010101010;
    r_input_signal[127] = 16'b0001011110111000;
    r_input_signal[128] = 16'b0001011011000011;
    r_input_signal[129] = 16'b0001010111001100;
    r_input_signal[130] = 16'b0001010011010011;
    r_input_signal[131] = 16'b0001001111010111;
    r_input_signal[132] = 16'b0001001011011000;
    r_input_signal[133] = 16'b0001000111011000;
    r_input_signal[134] = 16'b0001000011010110;
    r_input_signal[135] = 16'b0000111111010010;
    r_input_signal[136] = 16'b0000111011001100;
    r_input_signal[137] = 16'b0000110111000100;
    r_input_signal[138] = 16'b0000110010111011;
    r_input_signal[139] = 16'b0000101110110000;
    r_input_signal[140] = 16'b0000101010100101;
    r_input_signal[141] = 16'b0000100110010111;
    r_input_signal[142] = 16'b0000100010001001;
    r_input_signal[143] = 16'b0000011101111010;
    r_input_signal[144] = 16'b0000011001101010;
    r_input_signal[145] = 16'b0000010101011010;
    r_input_signal[146] = 16'b0000010001001000;
    r_input_signal[147] = 16'b0000001100110110;
    r_input_signal[148] = 16'b0000001000100100;
    r_input_signal[149] = 16'b0000000100010010;
    r_input_signal[150] = 16'b0000000000000000;
    r_input_signal[151] = 16'b1111111011101110;
    r_input_signal[152] = 16'b1111110111011100;
    r_input_signal[153] = 16'b1111110011001010;
    r_input_signal[154] = 16'b1111101110111000;
    r_input_signal[155] = 16'b1111101010100110;
    r_input_signal[156] = 16'b1111100110010110;
    r_input_signal[157] = 16'b1111100010000110;
    r_input_signal[158] = 16'b1111011101110111;
    r_input_signal[159] = 16'b1111011001101001;
    r_input_signal[160] = 16'b1111010101011011;
    r_input_signal[161] = 16'b1111010001010000;
    r_input_signal[162] = 16'b1111001101000101;
    r_input_signal[163] = 16'b1111001000111100;
    r_input_signal[164] = 16'b1111000100110100;
    r_input_signal[165] = 16'b1111000000101110;
    r_input_signal[166] = 16'b1110111100101010;
    r_input_signal[167] = 16'b1110111000101000;
    r_input_signal[168] = 16'b1110110100101000;
    r_input_signal[169] = 16'b1110110000101001;
    r_input_signal[170] = 16'b1110101100101101;
    r_input_signal[171] = 16'b1110101000110100;
    r_input_signal[172] = 16'b1110100100111101;
    r_input_signal[173] = 16'b1110100001001000;
    r_input_signal[174] = 16'b1110011101010110;
    r_input_signal[175] = 16'b1110011001100111;
    r_input_signal[176] = 16'b1110010101111011;
    r_input_signal[177] = 16'b1110010010010010;
    r_input_signal[178] = 16'b1110001110101011;
    r_input_signal[179] = 16'b1110001011001000;
    r_input_signal[180] = 16'b1110000111101001;
    r_input_signal[181] = 16'b1110000100001100;
    r_input_signal[182] = 16'b1110000000110011;
    r_input_signal[183] = 16'b1101111101011110;
    r_input_signal[184] = 16'b1101111010001100;
    r_input_signal[185] = 16'b1101110110111110;
    r_input_signal[186] = 16'b1101110011110100;
    r_input_signal[187] = 16'b1101110000101110;
    r_input_signal[188] = 16'b1101101101101100;
    r_input_signal[189] = 16'b1101101010101110;
    r_input_signal[190] = 16'b1101100111110100;
    r_input_signal[191] = 16'b1101100100111111;
    r_input_signal[192] = 16'b1101100010001110;
    r_input_signal[193] = 16'b1101011111100001;
    r_input_signal[194] = 16'b1101011100111001;
    r_input_signal[195] = 16'b1101011010010101;
    r_input_signal[196] = 16'b1101010111110110;
    r_input_signal[197] = 16'b1101010101011100;
    r_input_signal[198] = 16'b1101010011000110;
    r_input_signal[199] = 16'b1101010000110101;
    r_input_signal[200] = 16'b1101001110101010;
    r_input_signal[201] = 16'b1101001100100011;
    r_input_signal[202] = 16'b1101001010100001;
    r_input_signal[203] = 16'b1101001000100101;
    r_input_signal[204] = 16'b1101000110101101;
    r_input_signal[205] = 16'b1101000100111011;
    r_input_signal[206] = 16'b1101000011001110;
    r_input_signal[207] = 16'b1101000001100110;
    r_input_signal[208] = 16'b1101000000000100;
    r_input_signal[209] = 16'b1100111110100111;
    r_input_signal[210] = 16'b1100111101001111;
    r_input_signal[211] = 16'b1100111011111101;
    r_input_signal[212] = 16'b1100111010110001;
    r_input_signal[213] = 16'b1100111001101001;
    r_input_signal[214] = 16'b1100111000101000;
    r_input_signal[215] = 16'b1100110111101100;
    r_input_signal[216] = 16'b1100110110110110;
    r_input_signal[217] = 16'b1100110110000101;
    r_input_signal[218] = 16'b1100110101011010;
    r_input_signal[219] = 16'b1100110100110101;
    r_input_signal[220] = 16'b1100110100010110;
    r_input_signal[221] = 16'b1100110011111100;
    r_input_signal[222] = 16'b1100110011101000;
    r_input_signal[223] = 16'b1100110011011001;
    r_input_signal[224] = 16'b1100110011010001;
    r_input_signal[225] = 16'b1100110011001110;
    r_input_signal[226] = 16'b1100110011010001;
    r_input_signal[227] = 16'b1100110011011001;
    r_input_signal[228] = 16'b1100110011101000;
    r_input_signal[229] = 16'b1100110011111100;
    r_input_signal[230] = 16'b1100110100010110;
    r_input_signal[231] = 16'b1100110100110101;
    r_input_signal[232] = 16'b1100110101011010;
    r_input_signal[233] = 16'b1100110110000101;
    r_input_signal[234] = 16'b1100110110110110;
    r_input_signal[235] = 16'b1100110111101100;
    r_input_signal[236] = 16'b1100111000101000;
    r_input_signal[237] = 16'b1100111001101001;
    r_input_signal[238] = 16'b1100111010110001;
    r_input_signal[239] = 16'b1100111011111101;
    r_input_signal[240] = 16'b1100111101001111;
    r_input_signal[241] = 16'b1100111110100111;
    r_input_signal[242] = 16'b1101000000000100;
    r_input_signal[243] = 16'b1101000001100110;
    r_input_signal[244] = 16'b1101000011001110;
    r_input_signal[245] = 16'b1101000100111011;
    r_input_signal[246] = 16'b1101000110101101;
    r_input_signal[247] = 16'b1101001000100101;
    r_input_signal[248] = 16'b1101001010100001;
    r_input_signal[249] = 16'b1101001100100011;
    r_input_signal[250] = 16'b1101001110101010;
    r_input_signal[251] = 16'b1101010000110101;
    r_input_signal[252] = 16'b1101010011000110;
    r_input_signal[253] = 16'b1101010101011100;
    r_input_signal[254] = 16'b1101010111110110;
    r_input_signal[255] = 16'b1101011010010101;
    r_input_signal[256] = 16'b1101011100111001;
    r_input_signal[257] = 16'b1101011111100001;
    r_input_signal[258] = 16'b1101100010001110;
    r_input_signal[259] = 16'b1101100100111111;
    r_input_signal[260] = 16'b1101100111110100;
    r_input_signal[261] = 16'b1101101010101110;
    r_input_signal[262] = 16'b1101101101101100;
    r_input_signal[263] = 16'b1101110000101110;
    r_input_signal[264] = 16'b1101110011110100;
    r_input_signal[265] = 16'b1101110110111110;
    r_input_signal[266] = 16'b1101111010001100;
    r_input_signal[267] = 16'b1101111101011110;
    r_input_signal[268] = 16'b1110000000110011;
    r_input_signal[269] = 16'b1110000100001100;
    r_input_signal[270] = 16'b1110000111101001;
    r_input_signal[271] = 16'b1110001011001000;
    r_input_signal[272] = 16'b1110001110101011;
    r_input_signal[273] = 16'b1110010010010010;
    r_input_signal[274] = 16'b1110010101111011;
    r_input_signal[275] = 16'b1110011001100111;
    r_input_signal[276] = 16'b1110011101010110;
    r_input_signal[277] = 16'b1110100001001000;
    r_input_signal[278] = 16'b1110100100111101;
    r_input_signal[279] = 16'b1110101000110100;
    r_input_signal[280] = 16'b1110101100101101;
    r_input_signal[281] = 16'b1110110000101001;
    r_input_signal[282] = 16'b1110110100101000;
    r_input_signal[283] = 16'b1110111000101000;
    r_input_signal[284] = 16'b1110111100101010;
    r_input_signal[285] = 16'b1111000000101110;
    r_input_signal[286] = 16'b1111000100110100;
    r_input_signal[287] = 16'b1111001000111100;
    r_input_signal[288] = 16'b1111001101000101;
    r_input_signal[289] = 16'b1111010001010000;
    r_input_signal[290] = 16'b1111010101011011;
    r_input_signal[291] = 16'b1111011001101001;
    r_input_signal[292] = 16'b1111011101110111;
    r_input_signal[293] = 16'b1111100010000110;
    r_input_signal[294] = 16'b1111100110010110;
    r_input_signal[295] = 16'b1111101010100110;
    r_input_signal[296] = 16'b1111101110111000;
    r_input_signal[297] = 16'b1111110011001010;
    r_input_signal[298] = 16'b1111110111011100;
    r_input_signal[299] = 16'b1111111011101110;    
    // 100 samples test
    // r_input_signal[0] = 16'b0000000000000000;
    // r_input_signal[1] = 16'b0000001100110110;
    // r_input_signal[2] = 16'b0000011001101010;
    // r_input_signal[3] = 16'b0000100110010111;
    // r_input_signal[4] = 16'b0000110010111011;
    // r_input_signal[5] = 16'b0000111111010010;
    // r_input_signal[6] = 16'b0001001011011000;
    // r_input_signal[7] = 16'b0001010111001100;
    // r_input_signal[8] = 16'b0001100010101010;
    // r_input_signal[9] = 16'b0001101101101110;
    // r_input_signal[10] = 16'b0001111000010111;
    // r_input_signal[11] = 16'b0010000010100010;
    // r_input_signal[12] = 16'b0010001100001100;
    // r_input_signal[13] = 16'b0010010101010010;
    // r_input_signal[14] = 16'b0010011101110010;
    // r_input_signal[15] = 16'b0010100101101011;
    // r_input_signal[16] = 16'b0010101100111010;
    // r_input_signal[17] = 16'b0010110011011101;
    // r_input_signal[18] = 16'b0010111001010011;
    // r_input_signal[19] = 16'b0010111110011010;
    // r_input_signal[20] = 16'b0011000010110001;
    // r_input_signal[21] = 16'b0011000110010111;
    // r_input_signal[22] = 16'b0011001001001010;
    // r_input_signal[23] = 16'b0011001011001011;
    // r_input_signal[24] = 16'b0011001100011000;
    // r_input_signal[25] = 16'b0011001100110010;
    // r_input_signal[26] = 16'b0011001100011000;
    // r_input_signal[27] = 16'b0011001011001011;
    // r_input_signal[28] = 16'b0011001001001010;
    // r_input_signal[29] = 16'b0011000110010111;
    // r_input_signal[30] = 16'b0011000010110001;
    // r_input_signal[31] = 16'b0010111110011010;
    // r_input_signal[32] = 16'b0010111001010011;
    // r_input_signal[33] = 16'b0010110011011101;
    // r_input_signal[34] = 16'b0010101100111010;
    // r_input_signal[35] = 16'b0010100101101011;
    // r_input_signal[36] = 16'b0010011101110010;
    // r_input_signal[37] = 16'b0010010101010010;
    // r_input_signal[38] = 16'b0010001100001100;
    // r_input_signal[39] = 16'b0010000010100010;
    // r_input_signal[40] = 16'b0001111000010111;
    // r_input_signal[41] = 16'b0001101101101110;
    // r_input_signal[42] = 16'b0001100010101010;
    // r_input_signal[43] = 16'b0001010111001100;
    // r_input_signal[44] = 16'b0001001011011000;
    // r_input_signal[45] = 16'b0000111111010010;
    // r_input_signal[46] = 16'b0000110010111011;
    // r_input_signal[47] = 16'b0000100110010111;
    // r_input_signal[48] = 16'b0000011001101010;
    // r_input_signal[49] = 16'b0000001100110110;
    // r_input_signal[50] = 16'b0000000000000000;
    // r_input_signal[51] = 16'b1111110011001010;
    // r_input_signal[52] = 16'b1111100110010110;
    // r_input_signal[53] = 16'b1111011001101001;
    // r_input_signal[54] = 16'b1111001101000101;
    // r_input_signal[55] = 16'b1111000000101110;
    // r_input_signal[56] = 16'b1110110100101000;
    // r_input_signal[57] = 16'b1110101000110100;
    // r_input_signal[58] = 16'b1110011101010110;
    // r_input_signal[59] = 16'b1110010010010010;
    // r_input_signal[60] = 16'b1110000111101001;
    // r_input_signal[61] = 16'b1101111101011110;
    // r_input_signal[62] = 16'b1101110011110100;
    // r_input_signal[63] = 16'b1101101010101110;
    // r_input_signal[64] = 16'b1101100010001110;
    // r_input_signal[65] = 16'b1101011010010101;
    // r_input_signal[66] = 16'b1101010011000110;
    // r_input_signal[67] = 16'b1101001100100011;
    // r_input_signal[68] = 16'b1101000110101101;
    // r_input_signal[69] = 16'b1101000001100110;
    // r_input_signal[70] = 16'b1100111101001111;
    // r_input_signal[71] = 16'b1100111001101001;
    // r_input_signal[72] = 16'b1100110110110110;
    // r_input_signal[73] = 16'b1100110100110101;
    // r_input_signal[74] = 16'b1100110011101000;
    // r_input_signal[75] = 16'b1100110011001110;
    // r_input_signal[76] = 16'b1100110011101000;
    // r_input_signal[77] = 16'b1100110100110101;
    // r_input_signal[78] = 16'b1100110110110110;
    // r_input_signal[79] = 16'b1100111001101001;
    // r_input_signal[80] = 16'b1100111101001111;
    // r_input_signal[81] = 16'b1101000001100110;
    // r_input_signal[82] = 16'b1101000110101101;
    // r_input_signal[83] = 16'b1101001100100011;
    // r_input_signal[84] = 16'b1101010011000110;
    // r_input_signal[85] = 16'b1101011010010101;
    // r_input_signal[86] = 16'b1101100010001110;
    // r_input_signal[87] = 16'b1101101010101110;
    // r_input_signal[88] = 16'b1101110011110100;
    // r_input_signal[89] = 16'b1101111101011110;
    // r_input_signal[90] = 16'b1110000111101001;
    // r_input_signal[91] = 16'b1110010010010010;
    // r_input_signal[92] = 16'b1110011101010110;
    // r_input_signal[93] = 16'b1110101000110100;
    // r_input_signal[94] = 16'b1110110100101000;
    // r_input_signal[95] = 16'b1111000000101110;
    // r_input_signal[96] = 16'b1111001101000101;
    // r_input_signal[97] = 16'b1111011001101001;
    // r_input_signal[98] = 16'b1111100110010110;
    // r_input_signal[99] = 16'b1111110011001010;
  end

  // device under test
  top_dsm_dac_order_1 #(
    .DATA_WIDTH(DATA_WIDTH)
  ) dut (
    .i_clk(r_clk),
    .i_rst_n(r_rst_n),
    .i_sample(r_sample),
    .i_data(r_data_in),
    .o_dac_out(w_bit_out)
  );

  always #5 r_clk = ~r_clk; // 100 MHz = 10ns period

  integer file;
  integer i;
  integer j;
  initial begin
    file = $fopen("bitstream.txt","w");
    r_rst_n = 0;
    r_data_in = 0;
    #20 r_rst_n = 1;

    for (i = 0; i < $size(r_input_signal); i = i + 1) begin
      for (j = 0; j < OSR; j = j + 1) begin
        r_data_in = r_input_signal[i];
        @(posedge r_clk);
        $fwrite(file, "%0d\n", w_bit_out);
      end
    end

    $fclose(file);
    $display("Done, bitstream written to bitstream.txt");
    $finish;
  end

endmodule