`timescale 1ns/1ps

module tb_dsm_order1 #(
  parameter integer DATA_WIDTH = 16
) (
  // reg clk = 0;
  // reg rst_n = 0;
  // reg [DATA_WIDTH-1:0] data_in;
  // wire bit_out
);

  localparam input_signal [15:0] =
  {
    "16'b0111111111111111",
    "16'b1000100000001000",
    "16'b1001000000001010",
    "16'b1001011111111011",
    "16'b1001111111010100",
    "16'b1010011110001101",
    "16'b1010111100011110",
    "16'b1011011001111111",
    "16'b1011110110101001",
    "16'b1100010010010101",
    "16'b1100101100111011",
    "16'b1101000110010110",
    "16'b1101011110011110",
    "16'b1101110101001101",
    "16'b1110001010011111",
    "16'b1110011110001100",
    "16'b1110110000010010",
    "16'b1111000000101001",
    "16'b1111001111010000",
    "16'b1111011100000001",
    "16'b1111100110111011",
    "16'b1111101111111001",
    "16'b1111110110111010",
    "16'b1111111011111100",
    "16'b1111111110111110",
    "16'b1111111111111111",
    "16'b1111111110111110",
    "16'b1111111011111100",
    "16'b1111110110111010",
    "16'b1111101111111001",
    "16'b1111100110111011",
    "16'b1111011100000001",
    "16'b1111001111010000",
    "16'b1111000000101001",
    "16'b1110110000010010",
    "16'b1110011110001100",
    "16'b1110001010011111",
    "16'b1101110101001101",
    "16'b1101011110011110",
    "16'b1101000110010110",
    "16'b1100101100111011",
    "16'b1100010010010101",
    "16'b1011110110101001",
    "16'b1011011001111111",
    "16'b1010111100011110",
    "16'b1010011110001101",
    "16'b1001111111010100",
    "16'b1001011111111011",
    "16'b1001000000001010",
    "16'b1000100000001000",
    "16'b0111111111111111",
    "16'b0111011111110110",
    "16'b0110111111110100",
    "16'b0110100000000011",
    "16'b0110000000101010",
    "16'b0101100001110001",
    "16'b0101000011100000",
    "16'b0100100101111111",
    "16'b0100001001010101",
    "16'b0011101101101001",
    "16'b0011010011000011",
    "16'b0010111001101000",
    "16'b0010100001100000",
    "16'b0010001010110001",
    "16'b0001110101011111",
    "16'b0001100001110010",
    "16'b0001001111101100",
    "16'b0000111111010101",
    "16'b0000110000101110",
    "16'b0000100011111101",
    "16'b0000011001000011",
    "16'b0000010000000101",
    "16'b0000001001000100",
    "16'b0000000100000010",
    "16'b0000000001000000",
    "16'b0000000000000000",
    "16'b0000000001000000",
    "16'b0000000100000010",
    "16'b0000001001000100",
    "16'b0000010000000101",
    "16'b0000011001000011",
    "16'b0000100011111101",
    "16'b0000110000101110",
    "16'b0000111111010101",
    "16'b0001001111101100",
    "16'b0001100001110010",
    "16'b0001110101011111",
    "16'b0010001010110001",
    "16'b0010100001100000",
    "16'b0010111001101000",
    "16'b0011010011000011",
    "16'b0011101101101001",
    "16'b0100001001010101",
    "16'b0100100101111111",
    "16'b0101000011100000",
    "16'b0101100001110001",
    "16'b0110000000101010",
    "16'b0110100000000011",
    "16'b0110111111110100",
    "16'b0111011111110110"
  };

  reg r_clk = 0;
  reg r_rst_n = 0;
  reg [DATA_WIDTH-1:0] r_data_in;
  wire w_bit_out;

  top_dsm_dac_older_1 #(.DATA_WIDTH(DATA_WIDTH)) dut (
    .i_clk(r_clk),
    .i_rst_n(r_rst_n),
    .i_data(r_data_in),
    .o_dac_out(w_bit_out)
  );

  // clock
  always #5 r_clk = ~r_clk; // 100 MHz = 10ns period

  integer file;
  initial begin
    file = $fopen("bitstream.txt","w");
    r_rst_n = 0;
    r_data_in = 0;
    #20 r_rst_n = 1;

    // DC test: feed a constant positive input (e.g., mid-scale)
    r_data_in = 4'sd3; // change to test different inputs
    repeat (1000) begin
      @(posedge r_clk);
      $fwrite(file, "%0d\n", w_bit_out);
    end

    $fclose(file);
    $display("Done, bitstream written to bitstream.txt");
    $finish;
  end
endmodule