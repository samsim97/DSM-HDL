`timescale 1ns/1ps

module tb_top_dsm_dac_order_1;

  parameter integer DATA_WIDTH = 8;
  localparam integer NUM_SAMPLES = 100;

  reg r_clk = 0;
  reg r_rst_n = 0;
  reg r_sample = 1;
  reg signed [DATA_WIDTH-1:0] r_data_in = 0;
  wire w_bit_out;

  reg signed [DATA_WIDTH-1:0] r_input_signal [0:NUM_SAMPLES-1];

  initial begin
    r_input_signal[0] = 16'b0000000000000000;
    r_input_signal[1] = 16'b0000001100110110;
    r_input_signal[2] = 16'b0000011001101010;
    r_input_signal[3] = 16'b0000100110010111;
    r_input_signal[4] = 16'b0000110010111011;
    r_input_signal[5] = 16'b0000111111010010;
    r_input_signal[6] = 16'b0001001011011000;
    r_input_signal[7] = 16'b0001010111001100;
    r_input_signal[8] = 16'b0001100010101010;
    r_input_signal[9] = 16'b0001101101101110;
    r_input_signal[10] = 16'b0001111000010111;
    r_input_signal[11] = 16'b0010000010100010;
    r_input_signal[12] = 16'b0010001100001100;
    r_input_signal[13] = 16'b0010010101010010;
    r_input_signal[14] = 16'b0010011101110010;
    r_input_signal[15] = 16'b0010100101101011;
    r_input_signal[16] = 16'b0010101100111010;
    r_input_signal[17] = 16'b0010110011011101;
    r_input_signal[18] = 16'b0010111001010011;
    r_input_signal[19] = 16'b0010111110011010;
    r_input_signal[20] = 16'b0011000010110001;
    r_input_signal[21] = 16'b0011000110010111;
    r_input_signal[22] = 16'b0011001001001010;
    r_input_signal[23] = 16'b0011001011001011;
    r_input_signal[24] = 16'b0011001100011000;
    r_input_signal[25] = 16'b0011001100110010;
    r_input_signal[26] = 16'b0011001100011000;
    r_input_signal[27] = 16'b0011001011001011;
    r_input_signal[28] = 16'b0011001001001010;
    r_input_signal[29] = 16'b0011000110010111;
    r_input_signal[30] = 16'b0011000010110001;
    r_input_signal[31] = 16'b0010111110011010;
    r_input_signal[32] = 16'b0010111001010011;
    r_input_signal[33] = 16'b0010110011011101;
    r_input_signal[34] = 16'b0010101100111010;
    r_input_signal[35] = 16'b0010100101101011;
    r_input_signal[36] = 16'b0010011101110010;
    r_input_signal[37] = 16'b0010010101010010;
    r_input_signal[38] = 16'b0010001100001100;
    r_input_signal[39] = 16'b0010000010100010;
    r_input_signal[40] = 16'b0001111000010111;
    r_input_signal[41] = 16'b0001101101101110;
    r_input_signal[42] = 16'b0001100010101010;
    r_input_signal[43] = 16'b0001010111001100;
    r_input_signal[44] = 16'b0001001011011000;
    r_input_signal[45] = 16'b0000111111010010;
    r_input_signal[46] = 16'b0000110010111011;
    r_input_signal[47] = 16'b0000100110010111;
    r_input_signal[48] = 16'b0000011001101010;
    r_input_signal[49] = 16'b0000001100110110;
    r_input_signal[50] = 16'b0000000000000000;
    r_input_signal[51] = 16'b1111110011001010;
    r_input_signal[52] = 16'b1111100110010110;
    r_input_signal[53] = 16'b1111011001101001;
    r_input_signal[54] = 16'b1111001101000101;
    r_input_signal[55] = 16'b1111000000101110;
    r_input_signal[56] = 16'b1110110100101000;
    r_input_signal[57] = 16'b1110101000110100;
    r_input_signal[58] = 16'b1110011101010110;
    r_input_signal[59] = 16'b1110010010010010;
    r_input_signal[60] = 16'b1110000111101001;
    r_input_signal[61] = 16'b1101111101011110;
    r_input_signal[62] = 16'b1101110011110100;
    r_input_signal[63] = 16'b1101101010101110;
    r_input_signal[64] = 16'b1101100010001110;
    r_input_signal[65] = 16'b1101011010010101;
    r_input_signal[66] = 16'b1101010011000110;
    r_input_signal[67] = 16'b1101001100100011;
    r_input_signal[68] = 16'b1101000110101101;
    r_input_signal[69] = 16'b1101000001100110;
    r_input_signal[70] = 16'b1100111101001111;
    r_input_signal[71] = 16'b1100111001101001;
    r_input_signal[72] = 16'b1100110110110110;
    r_input_signal[73] = 16'b1100110100110101;
    r_input_signal[74] = 16'b1100110011101000;
    r_input_signal[75] = 16'b1100110011001110;
    r_input_signal[76] = 16'b1100110011101000;
    r_input_signal[77] = 16'b1100110100110101;
    r_input_signal[78] = 16'b1100110110110110;
    r_input_signal[79] = 16'b1100111001101001;
    r_input_signal[80] = 16'b1100111101001111;
    r_input_signal[81] = 16'b1101000001100110;
    r_input_signal[82] = 16'b1101000110101101;
    r_input_signal[83] = 16'b1101001100100011;
    r_input_signal[84] = 16'b1101010011000110;
    r_input_signal[85] = 16'b1101011010010101;
    r_input_signal[86] = 16'b1101100010001110;
    r_input_signal[87] = 16'b1101101010101110;
    r_input_signal[88] = 16'b1101110011110100;
    r_input_signal[89] = 16'b1101111101011110;
    r_input_signal[90] = 16'b1110000111101001;
    r_input_signal[91] = 16'b1110010010010010;
    r_input_signal[92] = 16'b1110011101010110;
    r_input_signal[93] = 16'b1110101000110100;
    r_input_signal[94] = 16'b1110110100101000;
    r_input_signal[95] = 16'b1111000000101110;
    r_input_signal[96] = 16'b1111001101000101;
    r_input_signal[97] = 16'b1111011001101001;
    r_input_signal[98] = 16'b1111100110010110;
    r_input_signal[99] = 16'b1111110011001010;
  end

  // localparam input_signal [15:0] =
  // {
  //   "16'b0111111111111111",
  //   "16'b1000100000001000",
  //   "16'b1001000000001010",
  //   "16'b1001011111111011",
  //   "16'b1001111111010100",
  //   "16'b1010011110001101",
  //   "16'b1010111100011110",
  //   "16'b1011011001111111",
  //   "16'b1011110110101001",
  //   "16'b1100010010010101",
  //   "16'b1100101100111011",
  //   "16'b1101000110010110",
  //   "16'b1101011110011110",
  //   "16'b1101110101001101",
  //   "16'b1110001010011111",
  //   "16'b1110011110001100",
  //   "16'b1110110000010010",
  //   "16'b1111000000101001",
  //   "16'b1111001111010000",
  //   "16'b1111011100000001",
  //   "16'b1111100110111011",
  //   "16'b1111101111111001",
  //   "16'b1111110110111010",
  //   "16'b1111111011111100",
  //   "16'b1111111110111110",
  //   "16'b1111111111111111",
  //   "16'b1111111110111110",
  //   "16'b1111111011111100",
  //   "16'b1111110110111010",
  //   "16'b1111101111111001",
  //   "16'b1111100110111011",
  //   "16'b1111011100000001",
  //   "16'b1111001111010000",
  //   "16'b1111000000101001",
  //   "16'b1110110000010010",
  //   "16'b1110011110001100",
  //   "16'b1110001010011111",
  //   "16'b1101110101001101",
  //   "16'b1101011110011110",
  //   "16'b1101000110010110",
  //   "16'b1100101100111011",
  //   "16'b1100010010010101",
  //   "16'b1011110110101001",
  //   "16'b1011011001111111",
  //   "16'b1010111100011110",
  //   "16'b1010011110001101",
  //   "16'b1001111111010100",
  //   "16'b1001011111111011",
  //   "16'b1001000000001010",
  //   "16'b1000100000001000",
  //   "16'b0111111111111111",
  //   "16'b0111011111110110",
  //   "16'b0110111111110100",
  //   "16'b0110100000000011",
  //   "16'b0110000000101010",
  //   "16'b0101100001110001",
  //   "16'b0101000011100000",
  //   "16'b0100100101111111",
  //   "16'b0100001001010101",
  //   "16'b0011101101101001",
  //   "16'b0011010011000011",
  //   "16'b0010111001101000",
  //   "16'b0010100001100000",
  //   "16'b0010001010110001",
  //   "16'b0001110101011111",
  //   "16'b0001100001110010",
  //   "16'b0001001111101100",
  //   "16'b0000111111010101",
  //   "16'b0000110000101110",
  //   "16'b0000100011111101",
  //   "16'b0000011001000011",
  //   "16'b0000010000000101",
  //   "16'b0000001001000100",
  //   "16'b0000000100000010",
  //   "16'b0000000001000000",
  //   "16'b0000000000000000",
  //   "16'b0000000001000000",
  //   "16'b0000000100000010",
  //   "16'b0000001001000100",
  //   "16'b0000010000000101",
  //   "16'b0000011001000011",
  //   "16'b0000100011111101",
  //   "16'b0000110000101110",
  //   "16'b0000111111010101",
  //   "16'b0001001111101100",
  //   "16'b0001100001110010",
  //   "16'b0001110101011111",
  //   "16'b0010001010110001",
  //   "16'b0010100001100000",
  //   "16'b0010111001101000",
  //   "16'b0011010011000011",
  //   "16'b0011101101101001",
  //   "16'b0100001001010101",
  //   "16'b0100100101111111",
  //   "16'b0101000011100000",
  //   "16'b0101100001110001",
  //   "16'b0110000000101010",
  //   "16'b0110100000000011",
  //   "16'b0110111111110100",
  //   "16'b0111011111110110"
  // };

  // device under test
  top_dsm_dac_older_1 #(
    .DATA_WIDTH(DATA_WIDTH)
  ) dut (
    .i_clk(r_clk),
    .i_rst_n(r_rst_n),
    .i_sample(r_sample),
    .i_data(r_data_in),
    .o_dac_out(w_bit_out)
  );

  always #5 r_clk = ~r_clk; // 100 MHz = 10ns period

  integer file;
  integer i;
  initial begin
    file = $fopen("bitstream.txt","w");
    r_rst_n = 0;
    r_data_in = 0;
    #20 r_rst_n = 1;

    for (i = 0; i < $size(r_input_signal); i = i + 1) begin
      r_data_in = r_input_signal[i];
      @(posedge r_clk);
      $fwrite(file, "%0d\n", w_bit_out);
    end

    $fclose(file);
    $display("Done, bitstream written to bitstream.txt");
    $finish;
  end

endmodule
// `timescale 1ns/1ps

// module tb_dsm_order1 #(
//   parameter integer DATA_WIDTH = 16
// ) (
//   // reg clk = 0;
//   // reg rst_n = 0;
//   // reg [DATA_WIDTH-1:0] data_in;
//   // wire bit_out
// );

//   localparam input_signal [15:0] =
//   {
//     "16'b0111111111111111",
//     "16'b1000100000001000",
//     "16'b1001000000001010",
//     "16'b1001011111111011",
//     "16'b1001111111010100",
//     "16'b1010011110001101",
//     "16'b1010111100011110",
//     "16'b1011011001111111",
//     "16'b1011110110101001",
//     "16'b1100010010010101",
//     "16'b1100101100111011",
//     "16'b1101000110010110",
//     "16'b1101011110011110",
//     "16'b1101110101001101",
//     "16'b1110001010011111",
//     "16'b1110011110001100",
//     "16'b1110110000010010",
//     "16'b1111000000101001",
//     "16'b1111001111010000",
//     "16'b1111011100000001",
//     "16'b1111100110111011",
//     "16'b1111101111111001",
//     "16'b1111110110111010",
//     "16'b1111111011111100",
//     "16'b1111111110111110",
//     "16'b1111111111111111",
//     "16'b1111111110111110",
//     "16'b1111111011111100",
//     "16'b1111110110111010",
//     "16'b1111101111111001",
//     "16'b1111100110111011",
//     "16'b1111011100000001",
//     "16'b1111001111010000",
//     "16'b1111000000101001",
//     "16'b1110110000010010",
//     "16'b1110011110001100",
//     "16'b1110001010011111",
//     "16'b1101110101001101",
//     "16'b1101011110011110",
//     "16'b1101000110010110",
//     "16'b1100101100111011",
//     "16'b1100010010010101",
//     "16'b1011110110101001",
//     "16'b1011011001111111",
//     "16'b1010111100011110",
//     "16'b1010011110001101",
//     "16'b1001111111010100",
//     "16'b1001011111111011",
//     "16'b1001000000001010",
//     "16'b1000100000001000",
//     "16'b0111111111111111",
//     "16'b0111011111110110",
//     "16'b0110111111110100",
//     "16'b0110100000000011",
//     "16'b0110000000101010",
//     "16'b0101100001110001",
//     "16'b0101000011100000",
//     "16'b0100100101111111",
//     "16'b0100001001010101",
//     "16'b0011101101101001",
//     "16'b0011010011000011",
//     "16'b0010111001101000",
//     "16'b0010100001100000",
//     "16'b0010001010110001",
//     "16'b0001110101011111",
//     "16'b0001100001110010",
//     "16'b0001001111101100",
//     "16'b0000111111010101",
//     "16'b0000110000101110",
//     "16'b0000100011111101",
//     "16'b0000011001000011",
//     "16'b0000010000000101",
//     "16'b0000001001000100",
//     "16'b0000000100000010",
//     "16'b0000000001000000",
//     "16'b0000000000000000",
//     "16'b0000000001000000",
//     "16'b0000000100000010",
//     "16'b0000001001000100",
//     "16'b0000010000000101",
//     "16'b0000011001000011",
//     "16'b0000100011111101",
//     "16'b0000110000101110",
//     "16'b0000111111010101",
//     "16'b0001001111101100",
//     "16'b0001100001110010",
//     "16'b0001110101011111",
//     "16'b0010001010110001",
//     "16'b0010100001100000",
//     "16'b0010111001101000",
//     "16'b0011010011000011",
//     "16'b0011101101101001",
//     "16'b0100001001010101",
//     "16'b0100100101111111",
//     "16'b0101000011100000",
//     "16'b0101100001110001",
//     "16'b0110000000101010",
//     "16'b0110100000000011",
//     "16'b0110111111110100",
//     "16'b0111011111110110"
//   };

//   reg r_clk = 0;
//   reg r_rst_n = 0;
//   reg [DATA_WIDTH-1:0] r_data_in;
//   wire w_bit_out;

//   top_dsm_dac_older_1 #(.DATA_WIDTH(DATA_WIDTH)) dut (
//     .i_clk(r_clk),
//     .i_rst_n(r_rst_n),
//     .i_data(r_data_in),
//     .o_dac_out(w_bit_out)
//   );

//   always #5 r_clk = ~r_clk; // 100 MHz = 10ns period

//   integer file;
//   integer i;
//   initial begin
//     file = $fopen("bitstream.txt","w");
//     r_rst_n = 0;
//     r_data_in = 0;
//     #20 r_rst_n = 1;

//     for (i = 0; i < $size(input_signal); i = i + 1) begin
//       r_data_in = input_signal[i];
//       @(posedge r_clk);
//       $fwrite(file, "%0d\n", w_bit_out);
//     end

//     $fclose(file);
//     $display("Done, bitstream written to bitstream.txt");
//     $finish;
//   end
// endmodule